----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 24.11.2017 12:45:41
-- Design Name: 
-- Module Name: audio_interface - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.package_dsed.all;
use IEEE.numeric_std.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity audio_interface is
Port (  clk_12megas : in STD_LOGIC;
        reset : in STD_LOGIC;
        --Recording ports
        --To/From the controller
        record_enable: in STD_LOGIC;
        sample_out: out STD_LOGIC_VECTOR (sample_size-1 downto 0);
        sample_out_ready: out STD_LOGIC;
        --To/From the microphone
        micro_clk : out STD_LOGIC;
        micro_data : in STD_LOGIC;
        micro_LR : out STD_LOGIC;
        --Playing ports
        --To/From the controller
        play_enable: in STD_LOGIC;
        sample_in: in std_logic_vector(sample_size-1 downto 0);
        sample_request: out std_logic;
        --To/From the mini-jack
        jack_sd : out STD_LOGIC;
        jack_pwm : out STD_LOGIC);
end audio_interface;


architecture Behavioral of audio_interface is

    component en_4_cycles is
    Port (  clk_12megas : in STD_LOGIC;
            reset : in STD_LOGIC;
            clk_3megas: out STD_LOGIC;
            en_2_cycles: out STD_LOGIC;
            en_4_cycles : out STD_LOGIC);
    end component;
    
    component FSMD_microphone is
        Port (  clk_12megas : in STD_LOGIC;
                reset : in STD_LOGIC;
                enable_4_cycles : in STD_LOGIC;
                micro_data : in STD_LOGIC;
                sample_out : out STD_LOGIC_VECTOR (sample_size-1 downto 0);
                sample_out_ready : out STD_LOGIC);
    end component;
    
    component pwm is
        port(
        clk_12megas: in std_logic;
        reset: in std_logic;
        en_2_cycles: in std_logic;
        sample_in: in std_logic_vector(sample_size-1 downto 0);
        sample_request: out std_logic;
        pwm_pulse: out std_logic
        );
    end component;
    
    signal enable_clk_3megas,enable_clk12megas_micro, enable_clk12megas_pwm, enable_2_cycles_in, enable_4_cycles_in, enable_2_cycles_out, enable_4_cycles_out: STD_LOGIC:='0';
    
begin

    en_4_c: en_4_cycles port map(
            clk_12megas=> clk_12megas,
            reset=> reset,
            clk_3megas => micro_clk, --enable_clk_3megas,
            en_2_cycles=> enable_2_cycles_in,
            en_4_cycles => enable_4_cycles_in
            );
    micro: FSMD_microphone port map(
            clk_12megas=> clk_12megas,
            reset=> reset,
            enable_4_cycles => enable_4_cycles_out,
            micro_data => micro_data,
            sample_out => sample_out,
            sample_out_ready => sample_out_ready
            );
    pwm_out: pwm port map(
            clk_12megas=> clk_12megas,
            reset=> reset,
            en_2_cycles=>enable_2_cycles_out,
            sample_in=>sample_in,
            sample_request=>sample_request,
            pwm_pulse => jack_pwm
            );
    
    jack_SD <='1';
    micro_LR <= '1';          
    enable_4_cycles_out <= enable_4_cycles_in and record_enable;
    enable_2_cycles_out <= enable_2_cycles_in and play_enable;
    
    
end Behavioral;
